* Full Adder SPICE Netlist
* Created: 04.Aug.2024 12:34:31

*.SCALE METER
*.GLOBAL vdd gnd

.SUBCKT Full_Adder VDD SUM Cout A B Cin GND
M37 n20 n25 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M38 n14 n20 n23 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M39 n23 n24 n14 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M66 n36 n13 n18 n3 C5NPMOS w=1.205e-6 l=3e-8 as=1.0845e-13 ps=2.77e-6 ad=1.62675e-13 pd=2.95e-6
M46 n17 n11 n5 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M58 n32 n21 n14 n0 C5NPMOS w=1.205e-6 l=3e-8 as=1.0845e-13 ps=2.77e-6 ad=1.62675e-13 pd=2.95e-6
M43 n26 n19 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M60 n11 n14 n12 n12 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M45 n10 n14 n18 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M71 n7 n27 n9 n9 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M48 n5 n13 n10 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M55 n20 n25 n28 n28 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M49 n5 n26 n17 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M61 n26 n19 n8 n8 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M53 n7 n27 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M50 n5 n20 n27 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M51 n10 n19 n5 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M41 n23 n25 n5 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M52 n15 n17 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M69 n3 n19 n36 n3 C5NPMOS w=1.205e-6 l=3e-8 as=1.0845e-13 ps=2.77e-6 ad=1.62675e-13 pd=2.95e-6
M40 n5 n21 n23 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M63 n18 n14 n33 n3 C5NPMOS w=1.205e-6 l=3e-8 as=1.0845e-13 ps=2.77e-6 ad=1.62675e-13 pd=2.95e-6
M47 n27 n29 n5 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M36 n21 n24 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M67 n17 n26 n34 n16 C5NPMOS w=1.2e-6 l=3e-8 as=8.4e-14 ps=2.68e-6 ad=1.8e-13 pd=3e-6
M59 n0 n25 n32 n0 C5NPMOS w=1.205e-6 l=3e-8 as=1.0845e-13 ps=2.77e-6 ad=1.62675e-13 pd=2.95e-6
M56 n31 n20 n0 n0 C5NPMOS w=1.205e-6 l=3e-8 as=1.0845e-13 ps=2.77e-6 ad=1.62675e-13 pd=2.95e-6
M65 n35 n29 n6 n6 C5NPMOS w=1.2e-6 l=3e-8 as=8.4e-14 ps=2.68e-6 ad=1.8e-13 pd=3e-6
M54 n21 n24 n1 n1 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M44 n18 n26 n10 n5 C5NNMOS w=2e-7 l=3e-8 as=1.4e-14 ps=6.8e-7 ad=3e-14 pd=1e-6
M62 n33 n26 n3 n3 C5NPMOS w=1.205e-6 l=3e-8 as=1.0845e-13 ps=2.77e-6 ad=1.62675e-13 pd=2.95e-6
M70 n15 n17 n2 n2 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M57 n14 n24 n31 n0 C5NPMOS w=1.205e-6 l=3e-8 as=1.0845e-13 ps=2.77e-6 ad=1.62675e-13 pd=2.95e-6
M68 n27 n20 n35 n6 C5NPMOS w=1.2e-6 l=3e-8 as=8.4e-14 ps=2.68e-6 ad=1.8e-13 pd=3e-6
M42 n11 n14 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M64 n34 n11 n16 n16 C5NPMOS w=1.2e-6 l=3e-8 as=8.4e-14 ps=2.68e-6 ad=1.8e-13 pd=3e-6
.ENDS Full_Adder

* Top-level netlist
VDD VDD 0 DC 5
GND GND 0 DC 0
VIN_A A 0 PULSE(0 5 0 1n 1n 10n 20n)
VIN_B B 0 PULSE(0 5 0 1n 1n 10n 20n)
VIN_Cin Cin 0 PULSE(0 5 0 1n 1n 10n 20n)

XFA1 VDD SUM Cout A B Cin GND Full_Adder

* Simulation control
.TRAN 1n 100n
.END
