*******************************************************************************
* CDL netlist
*
* Library : Training
* Top Cell Name: Full Adder
* View Name: extracted
* Netlist created: 03.Aug.2024 15:30:53
*******************************************************************************

*.SCALE METER
*.GLOBAL vdd gnd

*******************************************************************************
* Library Name: Training
* Cell Name:    Full Adder
* View Name:    extracted
*******************************************************************************

.SUBCKT Full Adder

M37 n20 n25 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M38 n14 n20 n23 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M39 n23 n24 n14 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M66 n36 n13 n18 n3 C5NPMOS w=1.205e-6 l=3e-8 as=3.2535e-13 ps=2.95e-6 ad=2.169e-13 pd=2.77e-6
M46 n17 n11 n5 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M58 n32 n21 n14 n0 C5NPMOS w=1.205e-6 l=3e-8 as=3.2535e-13 ps=2.95e-6 ad=2.169e-13 pd=2.77e-6
M43 n26 n19 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M60 n11 n14 n12 n12 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M45 n10 n14 n18 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M71 n7 n27 n9 n9 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M48 n5 n13 n10 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M55 n20 n25 n28 n28 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M49 n5 n26 n17 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M61 n26 n19 n8 n8 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M53 n7 n27 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M50 n5 n20 n27 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M51 n10 n19 n5 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M41 n23 n25 n5 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M52 n15 n17 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M69 n3 n19 n36 n3 C5NPMOS w=1.205e-6 l=3e-8 as=3.2535e-13 ps=2.95e-6 ad=2.169e-13 pd=2.77e-6
M40 n5 n21 n23 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M63 n18 n14 n33 n3 C5NPMOS w=1.205e-6 l=3e-8 as=3.2535e-13 ps=2.95e-6 ad=2.169e-13 pd=2.77e-6
M47 n27 n29 n5 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M36 n21 n24 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M67 n17 n26 n34 n16 C5NPMOS w=1.2e-6 l=3e-8 as=3.6e-13 ps=3e-6 ad=1.68e-13 pd=2.68e-6
M59 n0 n25 n32 n0 C5NPMOS w=1.205e-6 l=3e-8 as=3.2535e-13 ps=2.95e-6 ad=2.169e-13 pd=2.77e-6
M56 n31 n20 n0 n0 C5NPMOS w=1.205e-6 l=3e-8 as=3.2535e-13 ps=2.95e-6 ad=2.169e-13 pd=2.77e-6
M65 n35 n29 n6 n6 C5NPMOS w=1.2e-6 l=3e-8 as=3.6e-13 ps=3e-6 ad=1.68e-13 pd=2.68e-6
M54 n21 n24 n1 n1 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M44 n18 n26 n10 n5 C5NNMOS w=2e-7 l=3e-8 as=5.4e-14 ps=9.4e-7 ad=3.5e-14 pd=7.5e-7
M62 n33 n26 n3 n3 C5NPMOS w=1.205e-6 l=3e-8 as=3.2535e-13 ps=2.95e-6 ad=2.169e-13 pd=2.77e-6
M70 n15 n17 n2 n2 C5NPMOS w=2.9e-7 l=3e-8 as=2.755e-14 ps=7.7e-7 ad=2.755e-14 pd=7.7e-7
M57 n14 n24 n31 n0 C5NPMOS w=1.205e-6 l=3e-8 as=3.2535e-13 ps=2.95e-6 ad=2.169e-13 pd=2.77e-6
M68 n27 n20 n35 n6 C5NPMOS w=1.2e-6 l=3e-8 as=3.6e-13 ps=3e-6 ad=1.68e-13 pd=2.68e-6
M42 n11 n14 n5 n5 C5NNMOS w=1.9e-7 l=3e-8 as=1.805e-14 ps=5.7e-7 ad=1.805e-14 pd=5.7e-7
M64 n34 n11 n16 n16 C5NPMOS w=1.2e-6 l=3e-8 as=3.6e-13 ps=3e-6 ad=1.68e-13 pd=2.68e-6
.ENDS
